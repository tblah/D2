// this calls all the individual tests


module Test();
    initial
    begin
        $display("Hello World");
    end

endmodule
