** Profile: "TESTBENCH-testsim"  [ \\ugsamba\tde1g14\D2\subtractor\teamg_orcad-PSpiceFiles\TESTBENCH\testsim.sim ] 

** Creating circuit file "testsim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "//ugsamba/tde1g14/D2/libraries/schematic/d2.lib" 
* From [PSPICE NETLIST] section of C:\Users\tde1g14\AppData\Local\Temp\16.6.0/PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ns 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\TESTBENCH.net" 


.END
